.INCLUDE /home/nmendez/asic/bag3_skywater130_workspace/skywater130/calibre_setup/source.added

*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM


* Copyright 2019-2021 SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* This code is *alternatively* available under a BSD-3-Clause license, see
* details in the README.md at the top level and the license text at
* https://github.com/google/skywater-pdk-libs-sky130_bag3_pr/blob/master/LICENSE.alternative
*
* SPDX-License-Identifier: BSD-3-Clause OR Apache 2.0

.SUBCKT nmos4_hv B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nhv l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_hvesd B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nhvesd l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_svt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_lvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nlowvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hv B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phv l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hvesd B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phvesd l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_svt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B pshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_lvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B plowvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phighvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B pshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT res_metal_1 MINUS PLUS
*.PININFO MINUS:B PLUS:B
RR0 PLUS MINUS mrm1  m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT res_metal_2 MINUS PLUS
*.PININFO MINUS:B PLUS:B
RR0 PLUS MINUS mrm2  m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT res_metal_3 MINUS PLUS
*.PININFO MINUS:B PLUS:B
RR0 PLUS MINUS mrm3  m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT res_metal_4 MINUS PLUS
*.PININFO MINUS:B PLUS:B
RR0 PLUS MINUS mrm4  m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT res_metal_5 MINUS PLUS
*.PININFO MINUS:B PLUS:B
RR0 PLUS MINUS mrm5  m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT res_standard BULK MINUS PLUS
*.PININFO BULK:B MINUS:B PLUS:B
xR0 PLUS MINUS BULK xhrpoly m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT res_high_res BULK MINUS PLUS
*.PININFO BULK:B MINUS:B PLUS:B
xR0 PLUS MINUS BULK xuhrpoly m=1 w=w*1.0e6 l=l*1.0e6
.ENDS

.SUBCKT mim_standard BOT TOP
*.PININFO BOT:B TOP:B
CC0 TOP BOT xcmimc2 w=unit_width*1.0e6 l=unit_height*1.0e6 m=num_rows*num_cols
.ENDS

.SUBCKT mim_45 BOT TOP
*.PININFO BOT:B TOP:B
CC0 TOP BOT xcmimc2 w=unit_width*1.0e6 l=unit_height*1.0e6 m=num_rows*num_cols
.ENDS

.SUBCKT mim_34 BOT TOP
*.PININFO BOT:B TOP:B
CC0 TOP BOT xcmimc1 w=unit_width*1.0e6 l=unit_height*1.0e6 m=num_rows*num_cols
.ENDS


.SUBCKT nmos4_standard_w84_l30_seg4 b d g s
*.PININFO b:B d:B g:B s:B
XN b d g s / nmos4_standard l=150n nf=4 w=420n
.ENDS


.SUBCKT pmos4_standard_w110_l30_seg4 b d g s
*.PININFO b:B d:B g:B s:B
XP b d g s / pmos4_standard l=150n nf=4 w=550n
.ENDS


.SUBCKT inv in out VDD VSS
*.PININFO in:I out:O VDD:B VSS:B
XN VSS out in VSS / nmos4_standard_w84_l30_seg4
XP VDD out in VDD / pmos4_standard_w110_l30_seg4
.ENDS


.SUBCKT nmos4_standard_w84_l30_seg8 b d g s
*.PININFO b:B d:B g:B s:B
XN b d g s / nmos4_standard l=150n nf=8 w=420n
.ENDS


.SUBCKT pmos4_standard_w110_l30_seg8 b d g s
*.PININFO b:B d:B g:B s:B
XP b d g s / pmos4_standard l=150n nf=8 w=550n
.ENDS


.SUBCKT inv_1 in out VDD VSS
*.PININFO in:I out:O VDD:B VSS:B
XN VSS out in VSS / nmos4_standard_w84_l30_seg8
XP VDD out in VDD / pmos4_standard_w110_l30_seg8
.ENDS


.SUBCKT AA_inv_chain in out outb VDD VSS
*.PININFO in:I out:O outb:O VDD:B VSS:B
XINV0 in outb VDD VSS / inv
XINV1 outb out VDD VSS / inv_1
.ENDS
